module ExtendLoad
	(input logic [63:0] Ent_mem,
	 input logic [2:0] Seletor,
	 output logic [63:0] Saida);
	

	always_comb begin
		case(Seletor)
			// LD
			3'd0: begin
				Saida[63]=Ent_mem[63];
				Saida[62]=Ent_mem[62];
				Saida[61]=Ent_mem[61];
				Saida[60]=Ent_mem[60];
				Saida[59]=Ent_mem[59];
				Saida[58]=Ent_mem[58];
				Saida[57]=Ent_mem[57];
				Saida[56]=Ent_mem[56];
				Saida[55]=Ent_mem[55];
				Saida[54]=Ent_mem[54];
				Saida[53]=Ent_mem[53];
				Saida[52]=Ent_mem[52];
				Saida[51]=Ent_mem[51];
				Saida[50]=Ent_mem[50];
				Saida[49]=Ent_mem[49];
				Saida[48]=Ent_mem[48];
				Saida[47]=Ent_mem[47];
				Saida[46]=Ent_mem[46];
				Saida[45]=Ent_mem[45];
				Saida[44]=Ent_mem[44];
				Saida[43]=Ent_mem[43];
				Saida[42]=Ent_mem[42];
				Saida[41]=Ent_mem[41];
				Saida[40]=Ent_mem[40];
				Saida[39]=Ent_mem[39];
				Saida[38]=Ent_mem[38];
				Saida[37]=Ent_mem[37];
				Saida[36]=Ent_mem[36];
				Saida[35]=Ent_mem[35];
				Saida[34]=Ent_mem[34];
				Saida[33]=Ent_mem[33];
				Saida[32]=Ent_mem[32];
				Saida[31]=Ent_mem[31];
				Saida[30]=Ent_mem[30];
				Saida[29]=Ent_mem[29];
				Saida[28]=Ent_mem[28];
				Saida[27]=Ent_mem[27];
				Saida[26]=Ent_mem[26];
				Saida[25]=Ent_mem[25];
				Saida[24]=Ent_mem[24];
				Saida[23]=Ent_mem[23];
				Saida[22]=Ent_mem[22];
				Saida[21]=Ent_mem[21];
				Saida[20]=Ent_mem[20];
				Saida[19]=Ent_mem[19];
				Saida[18]=Ent_mem[18];
				Saida[17]=Ent_mem[17];
				Saida[16]=Ent_mem[16];
				Saida[15]=Ent_mem[15];
				Saida[14]=Ent_mem[14];
				Saida[13]=Ent_mem[13];
				Saida[12]=Ent_mem[12];
				Saida[11]=Ent_mem[11];
				Saida[10]=Ent_mem[10];
				Saida[9]=Ent_mem[9];
				Saida[8]=Ent_mem[8];
				Saida[7]=Ent_mem[7];
				Saida[6]=Ent_mem[6];
				Saida[5]=Ent_mem[5];
				Saida[4]=Ent_mem[4];
				Saida[3]=Ent_mem[3];
				Saida[2]=Ent_mem[2];
				Saida[1]=Ent_mem[1];
				Saida[0]=Ent_mem[0];
			end

			// LW
			3'd1: begin
				Saida[63]=Ent_mem[31];
				Saida[62]=Ent_mem[31];
				Saida[61]=Ent_mem[31];
				Saida[60]=Ent_mem[31];
				Saida[59]=Ent_mem[31];
				Saida[58]=Ent_mem[31];
				Saida[57]=Ent_mem[31];
				Saida[56]=Ent_mem[31];
				Saida[55]=Ent_mem[31];
				Saida[54]=Ent_mem[31];
				Saida[53]=Ent_mem[31];
				Saida[52]=Ent_mem[31];
				Saida[51]=Ent_mem[31];
				Saida[50]=Ent_mem[31];
				Saida[49]=Ent_mem[31];
				Saida[48]=Ent_mem[31];
				Saida[47]=Ent_mem[31];
				Saida[46]=Ent_mem[31];
				Saida[45]=Ent_mem[31];
				Saida[44]=Ent_mem[31];
				Saida[43]=Ent_mem[31];
				Saida[42]=Ent_mem[31];
				Saida[41]=Ent_mem[31];
				Saida[40]=Ent_mem[31];
				Saida[39]=Ent_mem[31];
				Saida[38]=Ent_mem[31];
				Saida[37]=Ent_mem[31];
				Saida[36]=Ent_mem[31];
				Saida[35]=Ent_mem[31];
				Saida[34]=Ent_mem[31];
				Saida[33]=Ent_mem[31];
				Saida[32]=Ent_mem[31];
				Saida[31]=Ent_mem[31];
				Saida[30]=Ent_mem[30];
				Saida[29]=Ent_mem[29];
				Saida[28]=Ent_mem[28];
				Saida[27]=Ent_mem[27];
				Saida[26]=Ent_mem[26];
				Saida[25]=Ent_mem[25];
				Saida[24]=Ent_mem[24];
				Saida[23]=Ent_mem[23];
				Saida[22]=Ent_mem[22];
				Saida[21]=Ent_mem[21];
				Saida[20]=Ent_mem[20];
				Saida[19]=Ent_mem[19];
				Saida[18]=Ent_mem[18];
				Saida[17]=Ent_mem[17];
				Saida[16]=Ent_mem[16];
				Saida[15]=Ent_mem[15];
				Saida[14]=Ent_mem[14];
				Saida[13]=Ent_mem[13];
				Saida[12]=Ent_mem[12];
				Saida[11]=Ent_mem[11];
				Saida[10]=Ent_mem[10];
				Saida[9]=Ent_mem[9];
				Saida[8]=Ent_mem[8];
				Saida[7]=Ent_mem[7];
				Saida[6]=Ent_mem[6];
				Saida[5]=Ent_mem[5];
				Saida[4]=Ent_mem[4];
				Saida[3]=Ent_mem[3];
				Saida[2]=Ent_mem[2];
				Saida[1]=Ent_mem[1];
				Saida[0]=Ent_mem[0];
			end

			// LH
	        	3'd2: begin
				Saida[63]=Ent_mem[15];
				Saida[62]=Ent_mem[15];
				Saida[61]=Ent_mem[15];
				Saida[60]=Ent_mem[15];
				Saida[59]=Ent_mem[15];
				Saida[58]=Ent_mem[15];
				Saida[57]=Ent_mem[15];
				Saida[56]=Ent_mem[15];
				Saida[55]=Ent_mem[15];
				Saida[54]=Ent_mem[15];
				Saida[53]=Ent_mem[15];
				Saida[52]=Ent_mem[15];
				Saida[51]=Ent_mem[15];
				Saida[50]=Ent_mem[15];
				Saida[49]=Ent_mem[15];
				Saida[48]=Ent_mem[15];
				Saida[47]=Ent_mem[15];
				Saida[46]=Ent_mem[15];
				Saida[45]=Ent_mem[15];
				Saida[44]=Ent_mem[15];
				Saida[43]=Ent_mem[15];
				Saida[42]=Ent_mem[15];
				Saida[41]=Ent_mem[15];
				Saida[40]=Ent_mem[15];
				Saida[39]=Ent_mem[15];
				Saida[38]=Ent_mem[15];
				Saida[37]=Ent_mem[15];
				Saida[36]=Ent_mem[15];
				Saida[35]=Ent_mem[15];
				Saida[34]=Ent_mem[15];
				Saida[33]=Ent_mem[15];
				Saida[32]=Ent_mem[15];
				Saida[31]=Ent_mem[15];
				Saida[30]=Ent_mem[15];
				Saida[29]=Ent_mem[15];
				Saida[28]=Ent_mem[15];
				Saida[27]=Ent_mem[15];
				Saida[26]=Ent_mem[15];
				Saida[25]=Ent_mem[15];
				Saida[24]=Ent_mem[15];
				Saida[23]=Ent_mem[15];
				Saida[22]=Ent_mem[15];
				Saida[21]=Ent_mem[15];
				Saida[20]=Ent_mem[15];
				Saida[19]=Ent_mem[15];
				Saida[18]=Ent_mem[15];
				Saida[17]=Ent_mem[15];
				Saida[16]=Ent_mem[15];
				Saida[15]=Ent_mem[15];
				Saida[14]=Ent_mem[14];
				Saida[13]=Ent_mem[13];
				Saida[12]=Ent_mem[12];
				Saida[11]=Ent_mem[11];
				Saida[10]=Ent_mem[10];
				Saida[9]=Ent_mem[9];
				Saida[8]=Ent_mem[8];
				Saida[7]=Ent_mem[7];
				Saida[6]=Ent_mem[6];
				Saida[5]=Ent_mem[5];
				Saida[4]=Ent_mem[4];
				Saida[3]=Ent_mem[3];
				Saida[2]=Ent_mem[2];
				Saida[1]=Ent_mem[1];
				Saida[0]=Ent_mem[0];
			end

			// LB
		    3'd3: begin
				Saida[63]=Ent_mem[7];
				Saida[62]=Ent_mem[7];
				Saida[61]=Ent_mem[7];
				Saida[60]=Ent_mem[7];
				Saida[59]=Ent_mem[7];
				Saida[58]=Ent_mem[7];
				Saida[57]=Ent_mem[7];
				Saida[56]=Ent_mem[7];
				Saida[55]=Ent_mem[7];
				Saida[54]=Ent_mem[7];
				Saida[53]=Ent_mem[7];
				Saida[52]=Ent_mem[7];
				Saida[51]=Ent_mem[7];
				Saida[50]=Ent_mem[7];
				Saida[49]=Ent_mem[7];
				Saida[48]=Ent_mem[7];
				Saida[47]=Ent_mem[7];
				Saida[46]=Ent_mem[7];
				Saida[45]=Ent_mem[7];
				Saida[44]=Ent_mem[7];
				Saida[43]=Ent_mem[7];
				Saida[42]=Ent_mem[7];
				Saida[41]=Ent_mem[7];
				Saida[40]=Ent_mem[7];
				Saida[39]=Ent_mem[7];
				Saida[38]=Ent_mem[7];
				Saida[37]=Ent_mem[7];
				Saida[36]=Ent_mem[7];
				Saida[35]=Ent_mem[7];
				Saida[34]=Ent_mem[7];
				Saida[33]=Ent_mem[7];
				Saida[32]=Ent_mem[7];
				Saida[31]=Ent_mem[7];
				Saida[30]=Ent_mem[7];
				Saida[29]=Ent_mem[7];
				Saida[28]=Ent_mem[7];
				Saida[27]=Ent_mem[7];
				Saida[26]=Ent_mem[7];
				Saida[25]=Ent_mem[7];
				Saida[24]=Ent_mem[7];
				Saida[23]=Ent_mem[7];
				Saida[22]=Ent_mem[7];
				Saida[21]=Ent_mem[7];
				Saida[20]=Ent_mem[7];
				Saida[19]=Ent_mem[7];
				Saida[18]=Ent_mem[7];
				Saida[17]=Ent_mem[7];
				Saida[16]=Ent_mem[7];
				Saida[15]=Ent_mem[7];
				Saida[14]=Ent_mem[7];
				Saida[13]=Ent_mem[7];
				Saida[12]=Ent_mem[7];
				Saida[11]=Ent_mem[7];
				Saida[10]=Ent_mem[7];
				Saida[9]=Ent_mem[7];
				Saida[8]=Ent_mem[7];
				Saida[7]=Ent_mem[7];
				Saida[6]=Ent_mem[6];
				Saida[5]=Ent_mem[5];
				Saida[4]=Ent_mem[4];
				Saida[3]=Ent_mem[3];
				Saida[2]=Ent_mem[2];
				Saida[1]=Ent_mem[1];
				Saida[0]=Ent_mem[0];
			end

			// LWU
			3'd4: begin
				Saida[63]=0;
				Saida[62]=0;
				Saida[61]=0;
				Saida[60]=0;
				Saida[59]=0;
				Saida[58]=0;
				Saida[57]=0;
				Saida[56]=0;
				Saida[55]=0;
				Saida[54]=0;
				Saida[53]=0;
				Saida[52]=0;
				Saida[51]=0;
				Saida[50]=0;
				Saida[49]=0;
				Saida[48]=0;
				Saida[47]=0;
				Saida[46]=0;
				Saida[45]=0;
				Saida[44]=0;
				Saida[43]=0;
				Saida[42]=0;
				Saida[41]=0;
				Saida[40]=0;
				Saida[39]=0;
				Saida[38]=0;
				Saida[37]=0;
				Saida[36]=0;
				Saida[35]=0;
				Saida[34]=0;
				Saida[33]=0;
				Saida[32]=0;
				Saida[31]=Ent_mem[31];
				Saida[30]=Ent_mem[30];
				Saida[29]=Ent_mem[29];
				Saida[28]=Ent_mem[28];
				Saida[27]=Ent_mem[27];
				Saida[26]=Ent_mem[26];
				Saida[25]=Ent_mem[25];
				Saida[24]=Ent_mem[24];
				Saida[23]=Ent_mem[23];
				Saida[22]=Ent_mem[22];
				Saida[21]=Ent_mem[21];
				Saida[20]=Ent_mem[20];
				Saida[19]=Ent_mem[19];
				Saida[18]=Ent_mem[18];
				Saida[17]=Ent_mem[17];
				Saida[16]=Ent_mem[16];
				Saida[15]=Ent_mem[15];
				Saida[14]=Ent_mem[14];
				Saida[13]=Ent_mem[13];
				Saida[12]=Ent_mem[12];
				Saida[11]=Ent_mem[11];
				Saida[10]=Ent_mem[10];
				Saida[9]=Ent_mem[9];
				Saida[8]=Ent_mem[8];
				Saida[7]=Ent_mem[7];
				Saida[6]=Ent_mem[6];
				Saida[5]=Ent_mem[5];
				Saida[4]=Ent_mem[4];
				Saida[3]=Ent_mem[3];
				Saida[2]=Ent_mem[2];
				Saida[1]=Ent_mem[1];
				Saida[0]=Ent_mem[0];
			end

			// LHU
			3'd5: begin
				Saida[63]=0;
				Saida[62]=0;
				Saida[61]=0;
				Saida[60]=0;
				Saida[59]=0;
				Saida[58]=0;
				Saida[57]=0;
				Saida[56]=0;
				Saida[55]=0;
				Saida[54]=0;
				Saida[53]=0;
				Saida[52]=0;
				Saida[51]=0;
				Saida[50]=0;
				Saida[49]=0;
				Saida[48]=0;
				Saida[47]=0;
				Saida[46]=0;
				Saida[45]=0;
				Saida[44]=0;
				Saida[43]=0;
				Saida[42]=0;
				Saida[41]=0;
				Saida[40]=0;
				Saida[39]=0;
				Saida[38]=0;
				Saida[37]=0;
				Saida[36]=0;
				Saida[35]=0;
				Saida[34]=0;
				Saida[33]=0;
				Saida[32]=0;
				Saida[31]=0;
				Saida[30]=0;
				Saida[29]=0;
				Saida[28]=0;
				Saida[27]=0;
				Saida[26]=0;
				Saida[25]=0;
				Saida[24]=0;
				Saida[23]=0;
				Saida[22]=0;
				Saida[21]=0;
				Saida[20]=0;
				Saida[19]=0;
				Saida[18]=0;
				Saida[17]=0;
				Saida[16]=0;
				Saida[15]=Ent_mem[15];
				Saida[14]=Ent_mem[14];
				Saida[13]=Ent_mem[13];
				Saida[12]=Ent_mem[12];
				Saida[11]=Ent_mem[11];
				Saida[10]=Ent_mem[10];
				Saida[9]=Ent_mem[9];
				Saida[8]=Ent_mem[8];
				Saida[7]=Ent_mem[7];
				Saida[6]=Ent_mem[6];
				Saida[5]=Ent_mem[5];
				Saida[4]=Ent_mem[4];
				Saida[3]=Ent_mem[3];
				Saida[2]=Ent_mem[2];
				Saida[1]=Ent_mem[1];
				Saida[0]=Ent_mem[0];

			end

			// LBU
			3'd6: begin
				Saida[63]=0;
				Saida[62]=0;
				Saida[61]=0;
				Saida[60]=0;
				Saida[59]=0;
				Saida[58]=0;
				Saida[57]=0;
				Saida[56]=0;
				Saida[55]=0;
				Saida[54]=0;
				Saida[53]=0;
				Saida[52]=0;
				Saida[51]=0;
				Saida[50]=0;
				Saida[49]=0;
				Saida[48]=0;
				Saida[47]=0;
				Saida[46]=0;
				Saida[45]=0;
				Saida[44]=0;
				Saida[43]=0;
				Saida[42]=0;
				Saida[41]=0;
				Saida[40]=0;
				Saida[39]=0;
				Saida[38]=0;
				Saida[37]=0;
				Saida[36]=0;
				Saida[35]=0;
				Saida[34]=0;
				Saida[33]=0;
				Saida[32]=0;
				Saida[31]=0;
				Saida[30]=0;
				Saida[29]=0;
				Saida[28]=0;
				Saida[27]=0;
				Saida[26]=0;
				Saida[25]=0;
				Saida[24]=0;
				Saida[23]=0;
				Saida[22]=0;
				Saida[21]=0;
				Saida[20]=0;
				Saida[19]=0;
				Saida[18]=0;
				Saida[17]=0;
				Saida[16]=0;
				Saida[15]=0;
				Saida[14]=0;
				Saida[13]=0;
				Saida[12]=0;
				Saida[11]=0;
				Saida[10]=0;
				Saida[9]=0;
				Saida[8]=0;
				Saida[7]=Ent_mem[7];
				Saida[6]=Ent_mem[6];
				Saida[5]=Ent_mem[5];
				Saida[4]=Ent_mem[4];
				Saida[3]=Ent_mem[3];
				Saida[2]=Ent_mem[2];
				Saida[1]=Ent_mem[1];
				Saida[0]=Ent_mem[0];
			end
		endcase
	end
endmodule

module ExtendStore
	(input logic [63:0] Ent_mem,
	 input logic [63:0] Ent_alt,
	 input logic [1:0] Seletor,
	 output logic [63:0] Saida);
	

	always_comb begin
		case(Seletor)
			2'd0: begin
				Saida[63]=Ent_mem[63];
				Saida[62]=Ent_mem[62];
				Saida[61]=Ent_mem[61];
				Saida[60]=Ent_mem[60];
				Saida[59]=Ent_mem[59];
				Saida[58]=Ent_mem[58];
				Saida[57]=Ent_mem[57];
				Saida[56]=Ent_mem[56];
				Saida[55]=Ent_mem[55];
				Saida[54]=Ent_mem[54];
				Saida[53]=Ent_mem[53];
				Saida[52]=Ent_mem[52];
				Saida[51]=Ent_mem[51];
				Saida[50]=Ent_mem[50];
				Saida[49]=Ent_mem[49];
				Saida[48]=Ent_mem[48];
				Saida[47]=Ent_mem[47];
				Saida[46]=Ent_mem[46];
				Saida[45]=Ent_mem[45];
				Saida[44]=Ent_mem[44];
				Saida[43]=Ent_mem[43];
				Saida[42]=Ent_mem[42];
				Saida[41]=Ent_mem[41];
				Saida[40]=Ent_mem[40];
				Saida[39]=Ent_mem[39];
				Saida[38]=Ent_mem[38];
				Saida[37]=Ent_mem[37];
				Saida[36]=Ent_mem[36];
				Saida[35]=Ent_mem[35];
				Saida[34]=Ent_mem[34];
				Saida[33]=Ent_mem[33];
				Saida[32]=Ent_mem[32];
				Saida[31]=Ent_alt[31];
				Saida[30]=Ent_alt[30];
				Saida[29]=Ent_alt[29];
				Saida[28]=Ent_alt[28];
				Saida[27]=Ent_alt[27];
				Saida[26]=Ent_alt[26];
				Saida[25]=Ent_alt[25];
				Saida[24]=Ent_alt[24];
				Saida[23]=Ent_alt[23];
				Saida[22]=Ent_alt[22];
				Saida[21]=Ent_alt[21];
				Saida[20]=Ent_alt[20];
				Saida[19]=Ent_alt[19];
				Saida[18]=Ent_alt[18];
				Saida[17]=Ent_alt[17];
				Saida[16]=Ent_alt[16];
				Saida[15]=Ent_alt[15];
				Saida[14]=Ent_alt[14];
				Saida[13]=Ent_alt[13];
				Saida[12]=Ent_alt[12];
				Saida[11]=Ent_alt[11];
				Saida[10]=Ent_alt[10];
				Saida[9]=Ent_alt[9];
				Saida[8]=Ent_alt[8];
				Saida[7]=Ent_alt[7];
				Saida[6]=Ent_alt[6];
				Saida[5]=Ent_alt[5];
				Saida[4]=Ent_alt[4];
				Saida[3]=Ent_alt[3];
				Saida[2]=Ent_alt[2];
				Saida[1]=Ent_alt[1];
				Saida[0]=Ent_alt[0];
			end
		      2'd1: begin
				Saida[63]=Ent_mem[63];
				Saida[62]=Ent_mem[62];
				Saida[61]=Ent_mem[61];
				Saida[60]=Ent_mem[60];
				Saida[59]=Ent_mem[59];
				Saida[58]=Ent_mem[58];
				Saida[57]=Ent_mem[57];
				Saida[56]=Ent_mem[56];
				Saida[55]=Ent_mem[55];
				Saida[54]=Ent_mem[54];
				Saida[53]=Ent_mem[53];
				Saida[52]=Ent_mem[52];
				Saida[51]=Ent_mem[51];
				Saida[50]=Ent_mem[50];
				Saida[49]=Ent_mem[49];
				Saida[48]=Ent_mem[48];
				Saida[47]=Ent_mem[47];
				Saida[46]=Ent_mem[46];
				Saida[45]=Ent_mem[45];
				Saida[44]=Ent_mem[44];
				Saida[43]=Ent_mem[43];
				Saida[42]=Ent_mem[42];
				Saida[41]=Ent_mem[41];
				Saida[40]=Ent_mem[40];
				Saida[39]=Ent_mem[39];
				Saida[38]=Ent_mem[38];
				Saida[37]=Ent_mem[37];
				Saida[36]=Ent_mem[36];
				Saida[35]=Ent_mem[35];
				Saida[34]=Ent_mem[34];
				Saida[33]=Ent_mem[33];
				Saida[32]=Ent_mem[32];
				Saida[31]=Ent_mem[31];
				Saida[30]=Ent_mem[30];
				Saida[29]=Ent_mem[29];
				Saida[28]=Ent_mem[28];
				Saida[27]=Ent_mem[27];
				Saida[26]=Ent_mem[26];
				Saida[25]=Ent_mem[25];
				Saida[24]=Ent_mem[24];
				Saida[23]=Ent_mem[23];
				Saida[22]=Ent_mem[22];
				Saida[21]=Ent_mem[21];
				Saida[20]=Ent_mem[20];
				Saida[19]=Ent_mem[19];
				Saida[18]=Ent_mem[18];
				Saida[17]=Ent_mem[17];
				Saida[16]=Ent_mem[16];
				Saida[15]=Ent_alt[15];
				Saida[14]=Ent_alt[14];
				Saida[13]=Ent_alt[13];
				Saida[12]=Ent_alt[12];
				Saida[11]=Ent_alt[11];
				Saida[10]=Ent_alt[10];
				Saida[9]=Ent_alt[9];
				Saida[8]=Ent_alt[8];
				Saida[7]=Ent_alt[7];
				Saida[6]=Ent_alt[6];
				Saida[5]=Ent_alt[5];
				Saida[4]=Ent_alt[4];
				Saida[3]=Ent_alt[3];
				Saida[2]=Ent_alt[2];
				Saida[1]=Ent_alt[1];
				Saida[0]=Ent_alt[0];

			end
		    2'd2: begin
				Saida[63]=Ent_mem[63];
				Saida[62]=Ent_mem[62];
				Saida[61]=Ent_mem[61];
				Saida[60]=Ent_mem[60];
				Saida[59]=Ent_mem[59];
				Saida[58]=Ent_mem[58];
				Saida[57]=Ent_mem[57];
				Saida[56]=Ent_mem[56];
				Saida[55]=Ent_mem[55];
				Saida[54]=Ent_mem[54];
				Saida[53]=Ent_mem[53];
				Saida[52]=Ent_mem[52];
				Saida[51]=Ent_mem[51];
				Saida[50]=Ent_mem[50];
				Saida[49]=Ent_mem[49];
				Saida[48]=Ent_mem[48];
				Saida[47]=Ent_mem[47];
				Saida[46]=Ent_mem[46];
				Saida[45]=Ent_mem[45];
				Saida[44]=Ent_mem[44];
				Saida[43]=Ent_mem[43];
				Saida[42]=Ent_mem[42];
				Saida[41]=Ent_mem[41];
				Saida[40]=Ent_mem[40];
				Saida[39]=Ent_mem[39];
				Saida[38]=Ent_mem[38];
				Saida[37]=Ent_mem[37];
				Saida[36]=Ent_mem[36];
				Saida[35]=Ent_mem[35];
				Saida[34]=Ent_mem[34];
				Saida[33]=Ent_mem[33];
				Saida[32]=Ent_mem[32];
				Saida[31]=Ent_mem[31];
				Saida[30]=Ent_mem[30];
				Saida[29]=Ent_mem[29];
				Saida[28]=Ent_mem[28];
				Saida[27]=Ent_mem[27];
				Saida[26]=Ent_mem[26];
				Saida[25]=Ent_mem[25];
				Saida[24]=Ent_mem[24];
				Saida[23]=Ent_mem[23];
				Saida[22]=Ent_mem[22];
				Saida[21]=Ent_mem[21];
				Saida[20]=Ent_mem[20];
				Saida[19]=Ent_mem[19];
				Saida[18]=Ent_mem[18];
				Saida[17]=Ent_mem[17];
				Saida[16]=Ent_mem[16];
				Saida[15]=Ent_mem[15];
				Saida[14]=Ent_mem[14];
				Saida[13]=Ent_mem[13];
				Saida[12]=Ent_mem[12];
				Saida[11]=Ent_mem[11];
				Saida[10]=Ent_mem[10];
				Saida[9]=Ent_mem[9];
				Saida[8]=Ent_mem[8];	
				Saida[7]=Ent_alt[7];
				Saida[6]=Ent_alt[6];
				Saida[5]=Ent_alt[5];
				Saida[4]=Ent_alt[4];
				Saida[3]=Ent_alt[3];
				Saida[2]=Ent_alt[2];
				Saida[1]=Ent_alt[1];
				Saida[0]=Ent_alt[0];

			end
		endcase
	end
endmodule
